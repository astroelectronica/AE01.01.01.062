.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C1608C0G2A100D080AA_p.mod"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/FMMT597.spice.txt"
.include "models/SMAZ15.spice.txt"
.include "models/ZXCT1008.spice.txt"
XU2 /SN /PWR_IN /COCM ZXCT1008F
R3 /PWR_IN /PWR_OUT 0.04
R4 /PWR_IN /PWR_OUT 0.04
R7 /SN /PWR_OUT 10k
XU3 /PWR_IN /SN C1608C0G2A100D080AA_p
R1 /BASE 0 1.5Meg
R5 /FILTER 0 4.99k
R6 /FILTER 0 4.99k
R2 /OUT /FILTER 100
XU5 /OUT 0 C2012C0G2A102J060AA_p
Q1 /FILTER /BASE /COCM FMMT597
I1 /PWR_OUT 0 {ILOAD}
V1 /PWR_IN 0 {VIN}
XU1 /BASE /PWR_IN SMAZ15
XU4 0 /OUT DI_BZX84C4V7
.end
